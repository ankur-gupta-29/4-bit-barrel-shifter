module barrel_shifter(
  input wire [3:0] i,
  input wire [1:0] s,
  output reg [3:0] o
);


endmodule
